module AND(x,b,y);
    input [31:0] x,b;
    output [31:0] y;
    assign y=b&x;
endmodule
    