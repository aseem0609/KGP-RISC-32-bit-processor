module OR(a,b,x);
    input [31:0] a,b;
    output [31:0] x;
    assign x=a|b;
    
endmodule