module Memory(address,store,write_data,mem_out,reset,pc,IF,clk,gcd,instr,booth);
    input [31:0] address,write_data,pc;
    output [31:0] mem_out;
    output reg [31:0] IF;
    input store,clk,reset,gcd,instr,booth;
    reg [1023:0] mem;
    always @(posedge clk)begin
        if(reset) mem<=0;
        if(gcd)begin
            mem[31:0]<=32'b010000_00000_00001_00000_00000_000000;
            mem[63:32]<=32'b010000_00001_00001_00000_00000_000110;  //loads data to R1
            mem[95:64]<=32'b010000_00000_00010_00000_00000_000000;
            mem[127:96]<=32'b010000_00010_00010_00000_00000_001111; //loads data to r2
            mem[159:128]<=32'b110001_00000_00000_00000_00000_000000; 
            mem[191:160]<=32'b000000_00001_00010_00011_00000_000001;
            mem[223:192]<=32'b011010_00000_00011_00000_00001_100000;
            mem[255:224]<=32'b011100_00000_00011_00000_00010_100000;
            mem[287:256]<=32'b000000_00001_00010_00001_00000_000001;
            mem[319:288]<=32'b011001_00000_00000_11111_11101_100000;
            mem[351:320]<=32'b000000_00010_00001_00010_00000_000001;
            mem[383:352]<=32'b011001_00000_00000_11111_11100_100000;
            mem[415:384]<=32'b110001_00000_00000_00000_00000_000000;
            
            mem[447:416]<=32'b110000_00010_00000_00000_00000_000000;
        end
        if(booth)begin
            mem[31:0]<=32'b010000_00000_00001_00000_00000_000000;       //M
            mem[63:32]<=32'b010000_00001_00001_00000_00000_000110;
            mem[95:64]<=32'b010000_00000_00010_00000_00000_000000;
            mem[127:96]<=32'b010000_00010_00010_00000_00000_001111;     //Q
            mem[159:128]<=32'b010000_00000_00011_00000_00000_100000;    //move 32 to R3
            mem[191:160]<=32'b010000_00000_00100_00000_00000_000000;    //Q-1
            mem[223:192]<=32'b010000_00000_00101_00000_00000_000000;    //A
            mem[255:224]<=32'b010000_00000_01000_00000_000000_00000;    //move 0 to R8
            mem[287:256]<=32'b010000_01000_01000_00000_000000_00001;    //R8=1           
            mem[319:288]<=32'b000001_00000_01001_00000_01111_100000;    //LOAD R9,992(R0)(R9=mem[1023:992]={1'b1,31'b0})
            mem[351:320]<=32'b110001_00000_00000_00000_00000_000000;    //beginning of loop
            mem[383:352]<=32'b000000_00010_01000_00110_00000_000010;    //AND R6,R2,R8(Q0)
            mem[415:384]<=32'b011011_00000_00110_00000_00010_000000;    //if Q0>0,jump
            mem[447:416]<=32'b011011_00000_00100_00000_00000_100000;    //if Q-1>0,jump to A=A+M
            mem[479:448]<=32'b011001_00000_00000_00000_00010_100000;    //jump to arithmetic shift
            mem[511:480]<=32'b000000_00101_00001_00101_00000_000000;    //A=A+M
            mem[543:512]<=32'b011001_00000_00000_00000_00001_100000;    //jump to arithmetic shift
            mem[575:544]<=32'b011100_00000_00100_00000_00000_100000;    //if Q-1=0,jump to A=A-M
            mem[607:576]<=32'b011001_00000_00000_00000_00000_100000;    //jump to arithmetic shift
            mem[639:608]<=32'b000000_00101_00001_00101_00000_000001;    //A=A-M
            mem[671:640]<=32'b000000_00010_01000_00100_00000_000010;    //AND R4,R8,R2(Q-1=Q0)
            mem[703:672]<=32'b011000_00010_00010_00000_00000_000001;    //SRLI Q,#1
            mem[735:704]<=32'b000000_00101_01000_00111_00000_000010;    //AND R7,R5,R8(R7=A0)
            mem[767:736]<=32'b011100_00000_00111_00000_00000_100000;    //if R7=0,skip next command
            mem[799:768]<=32'b000000_00010_01001_00010_00000_000000;    //R2=R2+R9
            mem[831:800]<=32'b010111_00101_00101_00000_00000_000001;    //SRAI A,#1
            mem[863:832]<=32'b000000_00011_01000_00011_00000_000001;    //SUB R3,R3,R8(count--)
            mem[895:864]<=32'b011011_00000_00011_11111_10111_100000;    //if count>0,jump to start of loop
            mem[927:896]<=32'b110000_00010_00000_00000_00000_000000;    //halt
            mem[1023:992]<=32'b100000_00000_00000_00000_000000_00000;
        end
        if(store)begin
            mem[address+:32]<=write_data;
        end
        if(instr)IF<=mem[pc+:32];
    end
    assign mem_out=mem[address+:32];
endmodule
